VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NAND
  CLASS CORE ;
  FOREIGN NAND ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SITE unithd ;
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.310 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.175 2.105 0.345 2.635 ;
        RECT 2.415 2.105 2.585 2.635 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000 0.095 2.760 0.795 ;
        RECT 0.145 -0.085 0.315 0.095 ;
    END
  END VNB
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.175 0.085 0.345 0.615 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.480 1.300 0.880 1.650 ;
    END
  END A
  PIN B
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.470 1.040 1.900 1.350 ;
    END
  END B
  PIN X
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.663600 ;
    PORT
      LAYER li1 ;
        RECT 1.295 1.745 1.465 2.445 ;
        RECT 1.295 1.660 2.585 1.745 ;
        RECT 1.295 1.575 2.615 1.660 ;
        RECT 2.300 1.060 2.615 1.575 ;
        RECT 2.415 0.275 2.585 1.060 ;
    END
  END X
END NAND
END LIBRARY

