VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SIGN
  CLASS BLOCK ;
  FOREIGN SIGN ;
  ORIGIN 0.000 0.000 ;
  SIZE 736.000 BY 448.000 ;
  SITE unithd ;
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 2.450 4.000 5.550 444.000 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 730.450 4.000 733.550 444.000 ;
    END
  END vccd1
  OBS
      LAYER met1 ;
        RECT 48.000 368.000 176.000 400.000 ;
        RECT 48.000 272.000 80.000 304.000 ;
        RECT 112.000 272.000 144.000 368.000 ;
        RECT 48.000 240.000 144.000 272.000 ;
        RECT 208.000 336.000 240.000 400.000 ;
        RECT 304.000 336.000 336.000 400.000 ;
        RECT 208.000 304.000 336.000 336.000 ;
        RECT 208.000 240.000 240.000 304.000 ;
        RECT 304.000 240.000 336.000 304.000 ;
        RECT 400.000 272.000 432.000 400.000 ;
        RECT 448.000 272.000 480.000 336.000 ;
        RECT 496.000 272.000 528.000 400.000 ;
        RECT 400.000 256.000 528.000 272.000 ;
        RECT 560.000 368.000 688.000 400.000 ;
        RECT 560.000 272.000 592.000 368.000 ;
        RECT 624.000 304.000 688.000 336.000 ;
        RECT 656.000 272.000 688.000 304.000 ;
        RECT 416.000 240.000 512.000 256.000 ;
        RECT 560.000 240.000 688.000 272.000 ;
        RECT 48.000 176.000 176.000 208.000 ;
        RECT 48.000 80.000 80.000 176.000 ;
        RECT 112.000 112.000 176.000 144.000 ;
        RECT 144.000 80.000 176.000 112.000 ;
        RECT 48.000 48.000 176.000 80.000 ;
        RECT 208.000 80.000 240.000 208.000 ;
        RECT 400.000 176.000 528.000 208.000 ;
        RECT 560.000 192.000 656.000 208.000 ;
        RECT 560.000 176.000 688.000 192.000 ;
        RECT 400.000 80.000 432.000 176.000 ;
        RECT 560.000 144.000 592.000 176.000 ;
        RECT 656.000 144.000 688.000 176.000 ;
        RECT 560.000 112.000 688.000 144.000 ;
        RECT 560.000 80.000 592.000 112.000 ;
        RECT 656.000 80.000 688.000 112.000 ;
        RECT 208.000 48.000 336.000 80.000 ;
        RECT 400.000 48.000 528.000 80.000 ;
        RECT 560.000 64.000 688.000 80.000 ;
        RECT 560.000 48.000 656.000 64.000 ;
      LAYER met2 ;
        RECT 48.000 368.000 176.000 400.000 ;
        RECT 48.000 272.000 80.000 304.000 ;
        RECT 112.000 272.000 144.000 368.000 ;
        RECT 48.000 240.000 144.000 272.000 ;
        RECT 208.000 336.000 240.000 400.000 ;
        RECT 304.000 336.000 336.000 400.000 ;
        RECT 208.000 304.000 336.000 336.000 ;
        RECT 208.000 240.000 240.000 304.000 ;
        RECT 304.000 240.000 336.000 304.000 ;
        RECT 400.000 272.000 432.000 400.000 ;
        RECT 448.000 272.000 480.000 336.000 ;
        RECT 496.000 272.000 528.000 400.000 ;
        RECT 400.000 256.000 528.000 272.000 ;
        RECT 560.000 368.000 688.000 400.000 ;
        RECT 560.000 272.000 592.000 368.000 ;
        RECT 624.000 304.000 688.000 336.000 ;
        RECT 656.000 272.000 688.000 304.000 ;
        RECT 416.000 240.000 512.000 256.000 ;
        RECT 560.000 240.000 688.000 272.000 ;
        RECT 48.000 176.000 176.000 208.000 ;
        RECT 48.000 80.000 80.000 176.000 ;
        RECT 112.000 112.000 176.000 144.000 ;
        RECT 144.000 80.000 176.000 112.000 ;
        RECT 48.000 48.000 176.000 80.000 ;
        RECT 208.000 80.000 240.000 208.000 ;
        RECT 400.000 176.000 528.000 208.000 ;
        RECT 560.000 192.000 656.000 208.000 ;
        RECT 560.000 176.000 688.000 192.000 ;
        RECT 400.000 80.000 432.000 176.000 ;
        RECT 560.000 144.000 592.000 176.000 ;
        RECT 656.000 144.000 688.000 176.000 ;
        RECT 560.000 112.000 688.000 144.000 ;
        RECT 560.000 80.000 592.000 112.000 ;
        RECT 656.000 80.000 688.000 112.000 ;
        RECT 208.000 48.000 336.000 80.000 ;
        RECT 400.000 48.000 528.000 80.000 ;
        RECT 560.000 64.000 688.000 80.000 ;
        RECT 560.000 48.000 656.000 64.000 ;
      LAYER met3 ;
        RECT 48.000 368.000 176.000 400.000 ;
        RECT 48.000 272.000 80.000 304.000 ;
        RECT 112.000 272.000 144.000 368.000 ;
        RECT 48.000 240.000 144.000 272.000 ;
        RECT 208.000 336.000 240.000 400.000 ;
        RECT 304.000 336.000 336.000 400.000 ;
        RECT 208.000 304.000 336.000 336.000 ;
        RECT 208.000 240.000 240.000 304.000 ;
        RECT 304.000 240.000 336.000 304.000 ;
        RECT 400.000 272.000 432.000 400.000 ;
        RECT 448.000 272.000 480.000 336.000 ;
        RECT 496.000 272.000 528.000 400.000 ;
        RECT 400.000 256.000 528.000 272.000 ;
        RECT 560.000 368.000 688.000 400.000 ;
        RECT 560.000 272.000 592.000 368.000 ;
        RECT 624.000 304.000 688.000 336.000 ;
        RECT 656.000 272.000 688.000 304.000 ;
        RECT 416.000 240.000 512.000 256.000 ;
        RECT 560.000 240.000 688.000 272.000 ;
        RECT 48.000 176.000 176.000 208.000 ;
        RECT 48.000 80.000 80.000 176.000 ;
        RECT 112.000 112.000 176.000 144.000 ;
        RECT 144.000 80.000 176.000 112.000 ;
        RECT 48.000 48.000 176.000 80.000 ;
        RECT 208.000 80.000 240.000 208.000 ;
        RECT 400.000 176.000 528.000 208.000 ;
        RECT 560.000 192.000 656.000 208.000 ;
        RECT 560.000 176.000 688.000 192.000 ;
        RECT 400.000 80.000 432.000 176.000 ;
        RECT 560.000 144.000 592.000 176.000 ;
        RECT 656.000 144.000 688.000 176.000 ;
        RECT 560.000 112.000 688.000 144.000 ;
        RECT 560.000 80.000 592.000 112.000 ;
        RECT 656.000 80.000 688.000 112.000 ;
        RECT 208.000 48.000 336.000 80.000 ;
        RECT 400.000 48.000 528.000 80.000 ;
        RECT 560.000 64.000 688.000 80.000 ;
        RECT 560.000 48.000 656.000 64.000 ;
      LAYER met4 ;
        RECT 48.000 368.000 176.000 400.000 ;
        RECT 48.000 272.000 80.000 304.000 ;
        RECT 112.000 272.000 144.000 368.000 ;
        RECT 48.000 240.000 144.000 272.000 ;
        RECT 208.000 336.000 240.000 400.000 ;
        RECT 304.000 336.000 336.000 400.000 ;
        RECT 208.000 304.000 336.000 336.000 ;
        RECT 208.000 240.000 240.000 304.000 ;
        RECT 304.000 240.000 336.000 304.000 ;
        RECT 400.000 272.000 432.000 400.000 ;
        RECT 448.000 272.000 480.000 336.000 ;
        RECT 496.000 272.000 528.000 400.000 ;
        RECT 400.000 256.000 528.000 272.000 ;
        RECT 560.000 368.000 688.000 400.000 ;
        RECT 560.000 272.000 592.000 368.000 ;
        RECT 624.000 304.000 688.000 336.000 ;
        RECT 656.000 272.000 688.000 304.000 ;
        RECT 416.000 240.000 512.000 256.000 ;
        RECT 560.000 240.000 688.000 272.000 ;
        RECT 48.000 176.000 176.000 208.000 ;
        RECT 48.000 80.000 80.000 176.000 ;
        RECT 112.000 112.000 176.000 144.000 ;
        RECT 144.000 80.000 176.000 112.000 ;
        RECT 48.000 48.000 176.000 80.000 ;
        RECT 208.000 80.000 240.000 208.000 ;
        RECT 400.000 176.000 528.000 208.000 ;
        RECT 560.000 192.000 656.000 208.000 ;
        RECT 560.000 176.000 688.000 192.000 ;
        RECT 400.000 80.000 432.000 176.000 ;
        RECT 560.000 144.000 592.000 176.000 ;
        RECT 656.000 144.000 688.000 176.000 ;
        RECT 560.000 112.000 688.000 144.000 ;
        RECT 560.000 80.000 592.000 112.000 ;
        RECT 656.000 80.000 688.000 112.000 ;
        RECT 208.000 48.000 336.000 80.000 ;
        RECT 400.000 48.000 528.000 80.000 ;
        RECT 560.000 64.000 688.000 80.000 ;
        RECT 560.000 48.000 656.000 64.000 ;
  END
END SIGN
END LIBRARY

